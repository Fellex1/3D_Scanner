*****************************************************************
* SIEMENS SIPMOS Power Transistors                              *
* SPICE Library Version 1.0                                     *
*                                                               *
* Models provided by SIEMENS are not warranted by SIEMENS as    *
* fully representing all of the specifications and operating    *
* characteristics of the semiconductor product to which the     *
* model relates. The model describe the characteristics of a    * 
* typical device.                                               * 
* In all cases, the current data sheet information for a given  *
* device is the final design guideline and the only actual      *
* performance specification.                                    *
* Altough models can be a useful tool in evaluating device      *
* performance, they cannot model exact device performance under *
* all conditions, nor are they intended to replace bread-       *
* boarding for final verification. SIEMENS reserves the right   *
* to change models without prior notice.                        *
*                                                               *
* This library contains the following                           *
* SIEMENS SIPMOS Transistors:                                   *
*                                                               *
*  BUZ-342KL    BUZ-51       BUZ-71LGE    BUZ-74A               *
*               BUZ-91A      BUZ-72       BUZ-45B               *
*  BUZ-12       BUZ-92       BUZ-311      BUZ-72GE              *
*  BUZ-323      BUZ-344      BUZ-50B      BUZ-73AGE             *
*  BUZ-21       BUZ-100_1    BUZ-73       BUZ-173               *
*  BUZ-10       BUZ-61A      BUZ-345      BUZ-11GE              *
*  BUZ-40B      BUZ-76                    BUZ-100_2             *
*  BUZ-81       BUZ-356      BUZ-220      BUZ-101               *
*  BUZ-20       BUZ-22       BUZ-78       BUZ-102               *
*  BUZ-11_2     BUZ-30A      BUZ-10M      BUZ-342               *
*  BUZ-358      BUZ-325      BUZ-305      BUZ-104               *
*  BUZ-80A      BUZ-60       BUZ-272                            *
*  BUZ-84A      BUZ-326      BUZ-77A                            *
*  BUZ-171      BUZ-11       BUZ-341                            *
*  BUZ-41A      BUZ-346      BUZ-331                            *
*  BUZ-70       BUZ-53A      BUZ-350                            *
*  BUZ-71L      BUZ-271      BUZ-310                            *
*  BUZ-10L      BUZ-334      BUZ-31                             *
*  BUZ-64       BUZ-12AL     BUZ-90                             *
*  BUZ-71       BUZ-73L      BUZ-338                            *
*                                                               *
*                                                               *
*---------------------------------------------------------------*
* connections:    gate                                          *
*                 | source                                      *
*                 | | drain                                     *
*                 | | |                                         *
*.subckt BUZ-342  1 2 3                                         *
*---------------------------------------------------------------*
 
 
***********
*SRC=BUZ-342KL;BUZ-342KL;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-342KL 1 2 3
LS 5 2 7N
LD 97 3 5N
RG 95 96 7.4
RS 5 76 0.01
D342 76 97 DREV
.MODEL DREV D CJO=6N RS=20M TT=150N IS=300P BV=50
M342 98 96 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.883 KP=17.8
M2 96 98 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 98 96 8 8 MSW
COX 96 8 15N
DGD 8 98 DCGD
.MODEL DCGD D CJO=3.6N M=0.548 VJ=1.027
CGS 76 96 8N
RD 98 97 0.0038
LG 95 1 7N
.ENDS
*******
*SRC=BUZ-12;BUZ-12;MOSFETs N;Siemens;50V 42A 28mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-12 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 76 24M
D12 76 86 DREV
.MODEL DREV D CJO=2N RS=20M TT=1.8N IS=300P BV=50
M12 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.516 KP=39.13
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 4N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.9N M=0.556 VJ=1.131
CGS 76 11 1.77N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-323;BUZ-323;MOSFETs N;Siemens;400V 15A 0.3 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-323 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 18M
D323 76 95 DREV
.MODEL DREV D CJO=0.7N RS=20M TT=40N IS=300P BV=400
M323 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.398 KP=16.36
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.649N M=0.555 VJ=1.006
CGS 76 11 2N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-13.58 KP=0.314
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-21;BUZ-21;MOSFETs N;Siemens;100V 21A 85mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-21 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 52M
D21 76 95 DREV
.MODEL DREV D CJO=1.2N RS=20M TT=50N IS=300P BV=100
M21 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.644 KP=21.65
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2.8N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.092N M=0.571 VJ=1.058
CGS 76 11 1.2N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.52 KP=12.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-10;BUZ-10;MOSFETs N;Siemens;50V 23A 70mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-10 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 51M
D10 76 95 DREV
.MODEL DREV D CJO=0.65N RS=20M TT=2.2N IS=300P BV=50
M10 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.287 KP=19.15
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 0.5N
DGD 8 95 DCGD
.MODEL DCGD D CJO=0.5N M=0.513 VJ=1.098
CGS 76 11 0.7N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-40B;BUZ-40B;MOSFETs N;Siemens;500V 8.5A 0.8 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-40B 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 20M
D40B 76 95 DREV
.MODEL DREV D CJO=0.5N RS=20M TT=400N IS=300P BV=500
M40B 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.813 KP=5.282
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.05N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.421N M=0.579 VJ=1.038
CGS 76 11 1.8N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-15.87 KP=0.112
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-81;BUZ-81;MOSFETs N;Siemens;800V 4A 2.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-81 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 23M
D81 76 95 DREV
.MODEL DREV D CJO=0.4N RS=20M TT=625N IS=300P BV=800
M81 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.463 KP=3.263
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.265N M=0.495 VJ=0.975
CGS 76 11 1N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-24.99 KP=.022
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-20;BUZ-20;MOSFETs N;Siemens;100V 13.5A 0.2 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-20 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 77M
D20 76 95 DREV
.MODEL DREV D CJO=0.35N RS=20M TT=100N IS=300P BV=100
M20 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.515 KP=7.547
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.560N M=0.556 VJ=1.056
CGS 76 11 0.46N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.71 KP=4
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-11_2;BUZ-11_2;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-11_2 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 26M
D21L 76 95 DREV
.MODEL DREV D CJO=0.7N RS=20M TT=23N IS=300P BV=50
M21L 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.605 KP=26.6
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 0.86N
DGD 8 95 DCGD
.MODEL DCGD D CJO=0.862N M=0.52 VJ=1.037
CGS 76 11 0.85N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-358;BUZ-358;MOSFETs N;Siemens;1000V 4.5A 2.6 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-358 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 64M
D358 76 95 DREV
.MODEL DREV D CJO=0.27N RS=20M TT=800N IS=300P BV=1000
M358 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.587 KP=15.84
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.75N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.553N M=0.541 VJ=1.016
CGS 76 11 2N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-41.34 KP=0.016
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-80A;BUZ-80A;MOSFETs N;Siemens;800V 3A 3 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-80A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 3.9
RS 5 76 51M
D80A 76 95 DREV
.MODEL DREV D CJO=0.45N RS=20M TT=1000N IS=300P BV=800
M80A 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.525 KP=2.996
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 86 11 8 8 MSW
COX 11 8 2.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.171N M=0.545 VJ=1.022
CGS 76 11 1.55N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-26.5 KP=0.014
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-84A;BUZ-84A;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-84A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 17M
D84A 76 95 DREV
.MODEL DREV D CJO=0.35N RS=20M TT=700N IS=300P BV=800
M84A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.736 KP=5.583
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.1N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.668N M=0.556 VJ=1.019
CGS 76 11 1.76N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-33.83 KP=0.029
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-171;BUZ-171;MOSFETs P;Siemens;50V 8A 0.3 Ohm
*SYM=P-MOSFET
.SUBCKT BUZ-171 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 76 128M
D171 86 76 DREV
.MODEL DREV D CJO=1.5N RS=20M TT=29N IS=300P BV=50
M171 86 11 76 76 MBUZ
.MODEL MBUZ PMOS VTO=-3.245 KP=0.973
M2 11 86 8 8 MSW
.MODEL MSW PMOS VTO=-0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.313N
DGD 86 8 DCGD
.MODEL DCGD D CJO=1.313N M=0.521 VJ=0.7
CGS 76 11 0.85N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-41A;BUZ-41A;MOSFETs N;Siemens;500V 4.5A 1.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-41A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 31M
D41A 76 95 DREV
.MODEL DREV D CJO=0.28N RS=20M TT=500N IS=300P BV=500
M41A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.277 KP=7.765
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.6N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.209N M=0.564 VJ=1.035
CGS 76 11 0.79N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-17.57 KP=0.055
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-70;BUZ-70;MOSFETs N;Siemens;60V 12A 0.15 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-70 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 136M
D70 76 95 DREV
.MODEL DREV D CJO=0.4N RS=20M TT=8.3N IS=300P BV=60
M70 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.68 KP=13.67
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 0.7N
DGD 8 95 DCGD
.MODEL DCGD D CJO=0.213N M=0.45 VJ=1.03
CGS 76 11 0.35N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-71L;BUZ-71L;MOSFETs N;Siemens;50V 14A 0.1 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-71L 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 76 64M
D71L 76 86 DREV
.MODEL DREV D CJO=0.55N RS=20M TT=10.7N IS=300P BV=50
M71L 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=2.057 KP=26.47
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=1
M3 86 11 8 8 MSW
COX 11 8 0.15N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.373N M=0.484 VJ=1.048
CGS 76 11 0.55N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-10L;BUZ-10L;MOSFETs N;Siemens;50V 23A 70mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-10L 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 76 70M
D10L 76 86 DREV
.MODEL DREV D CJO=7N RS=20M TT=4N IS=300P BV=50
M10L 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=2.562 KP=1415
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 8N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.491N M=0.502 VJ=1.047
CGS 76 11 1.5N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-64;BUZ-64;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-64 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 30M
D64 76 95 DREV
.MODEL DREV D CJO=0.8N RS=20M TT=100N IS=300P BV=400
M64 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.737 KP=13.14
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.775N M=0.609 VJ=1.045
CGS 76 11 1.8N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-14.1 KP=0.27
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-71;BUZ-71;MOSFETs N;Siemens;50V 14A 0.1 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-71 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 90M
D71 76 95 DREV
.MODEL DREV D CJO=0.48N RS=20M TT=7.1N IS=300P BV=50
M71 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.354 KP=20.7
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 0.9N
DGD 8 95 DCGD
.MODEL DCGD D CJO=0.340N M=0.480 VJ=1.099
CGS 76 11 0.4N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-51;BUZ-51;MOSFETs N;Siemens;1000V 3.4A 4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-51 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 9.8
RS 5 76 1M
D51 76 95 DREV
.MODEL DREV D CJO=0.3N RS=20M TT=300N IS=300P BV=1000
M51 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.994 KP=1.859
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.3
M3 86 11 8 8 MSW
COX 11 8 0.8N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.268N M=0.537 VJ=1.014
CGS 76 11 1N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-40.65 KP=0.0075
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-91A;BUZ-91A;MOSFETs N;Siemens;600V 8A 0.9 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-91A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 18M
D91A 76 95 DREV
.MODEL DREV D CJO=0.6N RS=50M TT=500N IS=300P BV=600
M91A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.725 KP=6.555
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.458N M=0.579 VJ=1.035
CGS 76 11 1.48N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-21.84 KP=0.069
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-92;BUZ-92;MOSFETs N;Siemens;600V 3.3A 3 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-92 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 41M
D92 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=500N IS=300P BV=600
M92 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.875 KP=2.349
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.168N M=0.567 VJ=1.038
CGS 76 11 0.6N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-19.91 KP=0.027
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-344;BUZ-344;MOSFETs N;Siemens;600V 12A 0.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-344 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 22M
D344 76 95 DREV
.MODEL DREV D CJO=3N RS=20M TT=100N IS=300P BV=100
M344 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.36 KP=44.73
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 6N
DGD 8 86 DCGD
.MODEL DCGD D CJO=2.9N M=0.575 VJ=1.017
CGS 76 11 11N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-55.64 KP=3
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-100_1;BUZ-100_1;MOSFETs N;Siemens;50V 60A 18mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-100_1 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 95 14M
D100 95 86 DREV
.MODEL DREV D CJO=3N RS=20M TT=200N IS=300P BV=50
M100 76 11 95 95 MBUZ
.MODEL MBUZ NMOS VTO=3.85 KP=30.02
M2 11 76 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 76 11 8 8 MSW
COX 11 8 5N
DGD 8 76 DCGD
.MODEL DCGD D CJO=1.389N M=0.511 VJ=1.055
CGS 95 11 3.03N
MRDR 76 76 86 76 MVRD
.MODEL MVRD NMOS VTO=-84.79 KP=5.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-61A;BUZ-61A;MOSFETs N;Siemens;400V 11A 0.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-61A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 3M
D61A 76 95 DREV
.MODEL DREV D CJO=0.4N RS=20M TT=400N IS=300P BV=400
M61A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.748 KP=5.122
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.505N M=0.537 VJ=0.988
CGS 76 11 1.49N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-14.22 KP=0.20
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-76;BUZ-76;MOSFETs N;Siemens;400V 3A 1.8 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-76 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 98M
D76 76 95 DREV
.MODEL DREV D CJO=0.12N RS=20M TT=800N IS=300P BV=400
M76 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.51 KP=2.422
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 .33N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.136N M=0.497 VJ=0.982
CGS 76 11 0.48N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-14.63 KP=0.06
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-356;BUZ-356;MOSFETs N;Siemens;800V 5.3A 2 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-356 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 53M
D356 76 95 DREV
.MODEL DREV D CJO=0.55N RS=20M TT=300N IS=300P BV=800
M356 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.24 KP=6.863
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.365N M=0.48 VJ=0.96
CGS 76 11 4.3N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-25.73 KP=0.044
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-22;BUZ-22;MOSFETs N;Siemens;100V 34A 55mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-22 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 34M
D22 76 95 DREV
.MODEL DREV D CJO=0.7N RS=20M TT=10N IS=300P BV=100
M22 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.76 KP=16.39
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2.2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.264N M=0.52 VJ=0.991
CGS 76 11 1.27N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-16.44 KP=4.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-30A;BUZ-30A;MOSFETs N;Siemens;200V 21A 0.13 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-30A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 36M
D30A 76 95 DREV
.MODEL DREV D CJO=0.6N RS=20M TT=60N IS=300P BV=200
M30A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.316 KP=29.38
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.7N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.860N M=0.527 VJ=0.983
CGS 76 11 1.29N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-12.08 KP=1.4
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-325;BUZ-325;MOSFETs N;Siemens;400V 12.5A 0.35 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-325 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 24M
D325 76 95 DREV
.MODEL DREV D CJO=0.5N RS=20M TT=400N IS=300P BV=400
M30A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.232 KP=13.57
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.628N M=0.533 VJ=0.981
CGS 76 11 1.71N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-15.38 KP=0.25
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-60;BUZ-60;MOSFETs N;Siemens;400V 5.5A 1 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-60 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 19M
D60 76 95 DREV
.MODEL DREV D CJO=.25N RS=20M TT=900N IS=300P BV=400
M60 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.711 KP=3.721
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 .6N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.275N M=0.515 VJ=0.981
CGS 76 11 0.76N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-15.02 KP=0.107
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-326;BUZ-326;MOSFETs N;Siemens;400V 10.5A 0.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-326 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 24M
D326 76 95 DREV
.MODEL DREV D CJO=0.45N RS=20M TT=480N IS=300P BV=400
M326 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.329 KP=13.21
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.507N M=0.497 VJ=0.982
CGS 76 11 1.19N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-15.31 KP=0.23
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-11;BUZ-11;MOSFETs N;Siemens;50V 30A 40mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-11 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 76 22M
D11 76 86 DREV
.MODEL DREV D CJO=1.5N RS=20M TT=4.2N IS=300P BV=50
M11 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.315 KP=24.41
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 3N
DGD 8 95 DCGD
.MODEL DCGD D CJO=1.03N M=0.537 VJ=1.135
CGS 76 11 1.22N
M347 86 95 95 95 MVRD
.MODEL MVRD NMOS VTO=-15.6 KP=10.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-346;BUZ-346;MOSFETs N;Siemens;50V 58A 18mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-346 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 10M
D346 76 95 DREV
.MODEL DREV D CJO=5.2N RS=20M TT=5.2N IS=300P BV=50
M346 95 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.188 KP=86.71
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 13N
DGD 8 95 DCGD
.MODEL DCGD D CJO=3.25N M=0.61 VJ=1.054
CGS 76 11 4N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-53A;BUZ-53A;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-53A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 30M
D53A 76 95 DREV
.MODEL DREV D CJO=0.22N RS=20M TT=2000N IS=300P BV=1000
M53A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.294 KP=2.402
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.45N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.124N M=0.443 VJ=0.968
CGS 76 11 1.46N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-36.62 KP=0.007
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-271;BUZ-271;MOSFETs P;Siemens;50V 22A 0.15 Ohm
*SYM=P-MOSFET
.SUBCKT BUZ-271 1 2 3
LS 5 2 7N
LD 87 3 5N
RG 4 11 5.5M
RS 5 76 58M
D271 87 76 DREV
.MODEL DREV D CJO=2N RS=20M TT=200N IS=300P BV=50
M271 87 11 76 76 MBUZ
.MODEL MBUZ PMOS VTO=-3.1 KP=1.956
M2 11 87 8 8 MSW
.MODEL MSW PMOS VTO=-0.001 KP=5
M3 87 11 8 8 MSW
COX 11 8 4.3N
DGD 87 8 DCGD
.MODEL DCGD D CJO=4.659N M=0.855 VJ=1.046
CGS 76 11 2N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-334;BUZ-334;MOSFETs N;Siemens;600V 12A 0.5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-334 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 3M
D334 76 95 DREV
.MODEL DREV D CJO=1.2N RS=20M TT=500N IS=300P BV=600
M334 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.748 KP=6.535
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.826N M=0.604 VJ=1.014
CGS 76 11 3.02N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-23.94 KP=.098
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-12AL;BUZ-12AL;MOSFETs N;Siemens;50V 42A 35mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-12AL 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 7.4
RS 5 76 13M
D12AL 76 95 DREV
.MODEL DREV D CJO=2.5N RS=20M TT=20N IS=300P BV=50
M12AL 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=1.913 KP=73.81
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 86 11 8 8 MSW
COX 11 8 6N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.64N M=0.564 VJ=1.036
CGS 76 11 2.1N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-28.82 KP=6
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-73L;BUZ-73L;MOSFETs N;Siemens;200V 7A 0.4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-73L 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 6.3
RS 5 76 42M
D73L 76 95 DREV
.MODEL DREV D CJO=0.3N RS=20M TT=100N IS=300P BV=200
M73L 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=1.941 KP=10.94
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 86 11 8 8 MSW
COX 11 8 2.5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.371N M=0.57 VJ=1.036
CGS 76 11 0.6N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.66 KP=.465
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-71LGE;BUZ-71LGE;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-71LGE 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 9.3
RS 5 76 34M
D71L 76 95 DREV
.MODEL DREV D CJO=0.55N RS=20M TT=30N IS=300P BV=50
M71L 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=1.918 KP=15.59
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 86 11 8 8 MSW
COX 11 8 2.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.411N M=0.507 VJ=1.042
CGS 76 11 0.55N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-30.7 KP=1.1
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-72;BUZ-72;MOSFETs N;Siemens;100V 10A 0.2 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-72 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 96M
D72 76 95 DREV
.MODEL DREV D CJO=0.3N RS=20M TT=50N IS=300P BV=100
M72 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.716 KP=4.828
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.423N M=0.568 VJ=1.053
CGS 76 11 0.36N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-11.58 KP=1.3
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-311;BUZ-311;MOSFETs N;Siemens;1000V 2.5A 5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-311 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 91M
D311 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=2000N IS=300P BV=1000
M311 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.098 KP=3.683
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.35N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.115N M=0.438 VJ=0.968
CGS 76 11 1.5N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-65.26 KP=0.0034
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-50B;BUZ-50B;MOSFETs N;Siemens;1000V 2A 8 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-50B 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 107M
D50B 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=2000N IS=300P BV=1000
M50B 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.342 KP=4.093
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 86 11 8 8 MSW
COX 11 8 0.4N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.123N M=0.451 VJ=0.969
CGS 76 11 1.5N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-35.45 KP=0.0075
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-73;BUZ-73;MOSFETs N;Siemens;200V 7A 0.4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-73 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 75M
D73 76 95 DREV
.MODEL DREV D CJO=0.28N RS=20M TT=200N IS=300P BV=200
M73 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.308 KP=8.528
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.348N M=0.544 VJ=1.056
CGS 76 11 0.47N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-9.182 KP=0.59
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-345;BUZ-345;MOSFETs N;Siemens;100V 41A 45 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-345 1 2 3
LS 5 2 7N
LD 87 3 5N
RG 4 11 5.5M
RS 5 76 36M
D345 76 87 DREV
.MODEL DREV D CJO=1.2N RS=20M TT=4.5N IS=300P BV=100
M345 87 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.618 KP=31.3
M2 11 87 8 8 MSW
.MODEL MSW NMOS VTO=0.0005 KP=10
M3 87 11 8 8 MSW IC=300,0,0
COX 11 8 5.5N
DGD 8 87 DCGD
.MODEL DCGD D CJO=2.13N M=0.614 VJ=1.146
CGS 76 11 1.6N
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-220;BUZ-220;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-220 1 2 3
LS 5 2 7N
LD 71 3 5N
RG 4 11 5.5M
RS 5 76 43M
D220 76 71 DREV
.MODEL DREV D CJO=580P RS=20M TT=121N IS=300P BV=900
M220 87 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.517 KP=4.781
M2 11 87 8 8 MSW
.MODEL MSW NMOS VTO=0.0005 KP=5
M3 87 11 8 8 MSW
COX 11 8 3.8N
DGD 8 87 DCGD
.MODEL DCGD D CJO=580P M=0.62 VJ=1.131
CGS 76 11 4.1N
MDR 71 87 87 87 MVARD
.MODEL MVARD NMOS VTO=-27.07 KP=.038
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-78;BUZ-78;MOSFETs N;Siemens;800V 1.5A 8 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-78 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 9.8
RS 5 76 155M
D78 76 95 DREV
.MODEL DREV D CJO=0.1N RS=20M TT=500N IS=300P BV=800
M78 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.649 KP=2.584
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.4
M3 86 11 8 8 MSW
COX 11 8 1N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.123N M=0.54 VJ=1.02
CGS 76 11 0.34N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-28.66 KP=0.007
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-10M;BUZ-10M;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-10M 1 2 3
LS 5 2 7N
LD 97 3 5N
RG 95 96 17.9
RS 5 76 0.018
D10M 76 97 DREV
.MODEL DREV D CJO=0.7N RS=20M TT=150N IS=300P BV=50
M10M 98 96 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.864 KP=8.138
M2 96 98 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 98 96 8 8 MSW
COX 96 8 2N
DGD 8 98 DCGD
.MODEL DCGD D CJO=0.371N M=0.467 VJ=1.029
CGS 76 96 0.7N
RD 98 97 0.025
LG 95 1 7N
.ENDS
*******
*SRC=BUZ-305;BUZ-305;MOSFETs N;Siemens;800V 7.5A 1 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-305 1 2 3
LS 5 2 7N
LD 97 3 5N
RG 95 96 5.8
RS 5 76 0.044
D305 76 97 DREV
.MODEL DREV D CJO=0.75N RS=20M TT=150N IS=300P BV=800
M305 99 96 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.617 KP=10.163
M2 96 99 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.5
M3 99 96 8 8 MSW
COX 96 8 4N
DGD 8 99 DCGD
.MODEL DCGD D CJO=0.735N M=0.549 VJ=0.996
CGS 76 96 2.1N
MRDR 99 99 97 99 MVRD
.MODEL MVRD NMOS VTO=-53.44 KP=0.022
LG 95 1 7N
.ENDS
*******
*SRC=BUZ-272;BUZ-272;MOSFETs P;Siemens;100V 15A 0.3mOhm
*SYM=P-MOSFET
.SUBCKT BUZ-272 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 95 9.6
RS 5 76 56M
D272 86 76 DREV
.MODEL DREV D CJO=1.7N RS=20M TT=180N IS=300P BV=100
M272 102 95 76 76 MBUZ
.MODEL MBUZ PMOS VTO=-3.149 KP=1.761
M2 11 102 8 8 MSW
.MODEL MSW PMOS VTO=-0.001 KP=.5
M3 102 11 8 8 MSW
COX 11 8 700P
DGD 102 8 DCGD
.MODEL DCGD D CJO=692P M=0.659 VJ=1.029
CGS 76 95 2N
VGC 11 95 -10
* BESCHREIBT EINE IMPLANTIERTE LADUNG (VERSCHIEBT DIE EINSATZSPANNUNG)
MHELP 86 102 102 102 MVRD
.MODEL MVRD PMOS VTO=13 KP=0.8
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-77A;BUZ-77A;MOSFETs N;Siemens;600V 2.7A 4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-77A 1 2 3
LS 5 2 7N
LD 97 3 5N
RG 95 99 6.8
RS 5 76 0.029
D77A 76 97 DREV
.MODEL DREV D CJO=0.25N RS=20M TT=800N IS=300P BV=600
M77A 98 99 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.909 KP=1.283
M2 87 98 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.4
M3 98 87 8 8 MSW
COX 87 8 0.17N
DGD 8 98 DCGD
.MODEL DCGD D CJO=116.75P M=0.553 VJ=1.017
CGS 76 99 0.34N
VGC 87 99 3
MHELP 98 98 97 98 MVRD
.MODEL MVRD NMOS VTO=-21.01 KP=0.018
LG 95 1 7N
.ENDS
*******
*SRC=BUZ-341;BUZ-341;MOSFETs N;Siemens;200V 33A 70mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-341 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 14M
D341 76 95 DREV
.MODEL DREV D CJO=0.9N RS=20M TT=30N IS=300P BV=200
M341 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.248 KP=26.86
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2.7N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.547N M=0.522 VJ=0.977
CGS 76 11 2.5N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.85 KP=2.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-331;BUZ-331;MOSFETs N;Siemens;500V 8A 0.8 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-331 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 24M
D331 76 95 DREV
.MODEL DREV D CJO=0.4 RS=20M TT=600N IS=300P BV=500
M331 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.089 KP=9.144
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.353N M=0.498 VJ=0.983
CGS 76 11 1.24N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-17.9 KP=0.104
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-350;BUZ-350;MOSFETs N;Siemens;200V 22A 0.12 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-350 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 23M
D350 76 95 DREV
.MODEL DREV D CJO=.8N RS=20M TT=270N IS=300P BV=200
M350 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.366 KP=23.29
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=1.103N M=0.53 VJ=0.984
CGS 76 11 1.6N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.24 KP=1.65
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-310;BUZ-310;MOSFETs N;Siemens;1000V 2.5A 5 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-310 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 31M
D310 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=2000N IS=300P BV=1000
+
M310 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.118 KP=2.132
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.35N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.649N M=0.555 VJ=1.006
CGS 76 11 1.5N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-33.31 KP=0.007
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-31;BUZ-31;MOSFETs N;Siemens;200V 14.5A 0.2 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-31 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 28M
D31 76 95 DREV
.MODEL DREV D CJO=0.33N RS=20M TT=100N IS=300P BV=200
M31 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.048 KP=13.97
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.626N M=0.523 VJ=0.985
CGS 76 11 0.81N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-9.935 KP=1.08
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-90;BUZ-90;MOSFETs N;Siemens;600V 4.5A 1.6 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-90 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 20M
D90 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=750N IS=300P BV=600
M90 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.227 KP=4.485
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.5N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.197N M=0.48 VJ=0.977
CGS 76 11 0.7N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-24.69 KP=0.031
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-338;BUZ-338;MOSFETs N;Siemens;500V 13.5A 0.4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-338 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 14M
D338 76 95 DREV
.MODEL DREV D CJO=0.65N RS=20M TT=500N IS=300P BV=500
M338 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.53 KP=15.731
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.867N M=0.578 VJ=1.016
CGS 76 11 2.5N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-19.18 KP=0.175
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-74A;BUZ-74A;MOSFETs N;Siemens;500V 2.1A 4 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-74A 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 76M
D74A 76 95 DREV
.MODEL DREV D CJO=0.15N RS=20M TT=500N IS=300P BV=500
M74A 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.835 KP=1.768
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.38N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.136N M=0.534 VJ=1.014
CGS 76 11 0.47N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-18.14 KP=0.032
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-45B;BUZ-45B;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-45B 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 53M
D45B 76 95 DREV
.MODEL DREV D CJO=0.8N RS=20M TT=120N IS=300P BV=500
M45B 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.268 KP=9.404
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2.3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.753N M=0.575 VJ=1.046
CGS 76 11 4.15N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-18.48 KP=0.149
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-72GE;BUZ-72GE;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-72GE 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 96M
D72 76 95 DREV
.MODEL DREV D CJO=0.3N RS=20M TT=50N IS=300P BV=100
M72 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.716 KP=4.828
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.423N M=0.568 VJ=1.053
CGS 76 11 0.36N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-11.58 KP=1.3
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-73AGE;BUZ-73AGE;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-73AGE 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 60M
D73A 76 95 DREV
.MODEL DREV D CJO=0.2N RS=20M TT=100N IS=300P BV=200
M73 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=3.618 KP=3.398
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 1.2N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.279N M=0.60 VJ=0.965
CGS 76 11 0.36N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-10.05 KP=.33
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-173;BUZ-173;MOSFETs P;Siemens;200V 3.6A 1.5 Ohm
*SYM=P-MOSFET
.SUBCKT BUZ-173 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 95 5.5M
RS 5 76 129M
D173 86 76 DREV
.MODEL DREV D CJO=550P RS=20M TT=180N IS=300P BV=200
M173 102 95 76 76 MBUZ
.MODEL MBUZ PMOS VTO=-3.419 KP=0.986
M2 11 102 8 8 MSW
.MODEL MSW PMOS VTO=-0.001 KP=5
M3 102 11 8 8 MSW
COX 11 8 300P
DGD 102 8 DCGD
.MODEL DCGD D CJO=204P M=0.533 VJ=1.01
CGS 76 95 800P
VGC 11 95 -9
* BESCHREIBT EINE IMPLANTIERTE LADUNG (VERSCHIEBT DIE EINSATZSPANNUNG)
MHELP 86 102 102 102 MVRD
.MODEL MVRD PMOS VTO=14.79 KP=0.08
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-11GE;BUZ-11GE;MOSFETs N;Siemens;
*SYM=N-MOSFET
.SUBCKT BUZ-11GE 1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 16M
D11 76 95 DREV
.MODEL DREV D CJO=1.35N RS=20M TT=100N IS=300P BV=50
M11 86 11 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.38 KP=15.04
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 3N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.936N M=0.544 VJ=1.099
CGS 76 11 1.05N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-13.86 KP=8.8
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-100_2;BUZ-100_2;MOSFETs N;Siemens;50V 60A 18mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-100_2 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 96 2.292M
D100 96 86 DREV
.MODEL DREV D CJO=3N RS=20M TT=30N IS=300P BV=50
M100 95 11 96 96 MBUZ
.MODEL MBUZ NMOS VTO=3.496 KP=22.66
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 7.21N
DGD 8 95 DCGD
.MODEL DCGD D CJO=4.2962N M=0.5 VJ=1
CGS 96 11 2.7098N
MHELP 95 95 86 95 MVRD
.MODEL MVRD NMOS VTO=-3.875 KP=19.5
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-101;BUZ-101;MOSFETs N;Siemens;50V 29A 60mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-101 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 96 4.987M
D101 96 86 DREV
.MODEL DREV D CJO=0.70294N RS=20M TT=30N IS=300P BV=50
M101 95 11 96 96 MBUZ
.MODEL MBUZ NMOS VTO=3.394 KP=7.926
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 0.99N
DGD 8 95 DCGD
.MODEL DCGD D CJO=0.9904N M=0.5 VJ=1
CGS 96 11 0.62085N
MHELP 95 95 86 95 MVRD
.MODEL MVRD NMOS VTO=-2.6 KP=17.1
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-102;BUZ-102;MOSFETs N;Siemens;50V 42A 23mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-102 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 96 13.21M
D102 96 86 DREV
.MODEL DREV D CJO=2.06393N RS=20M TT=30N IS=300P BV=50
M102 95 11 96 96 MBUZ
.MODEL MBUZ NMOS VTO=3.123 KP=21.57
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 4.096N
DGD 8 95 DCGD
.MODEL DCGD D CJO=2.5964N M=0.5 VJ=1
CGS 96 11 1.53485N
MHELP 95 95 86 95 MVRD
.MODEL MVRD NMOS VTO=-7.776 KP=13
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-342;BUZ-342;MOSFETs N;Siemens;50V 60A 10mOhm
*SYM=N-MOSFET
.SUBCKT BUZ-342 1 2 3
LS 5 2 7N
LD 86 3 5N
RG 4 11 5.5M
RS 5 96 12.74M
D342 96 86 DREV
.MODEL DREV D CJO=7.49393N RS=20M TT=85N IS=300P BV=50
M342 95 11 96 96 MBUZ
.MODEL MBUZ NMOS VTO=4.137 KP=69.74
M2 11 95 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 95 11 8 8 MSW
COX 11 8 163.09N
DGD 8 95 DCGD
.MODEL DCGD D CJO=11.6664N M=0.5 VJ=1
CGS 96 11 7.23985N
MHELP 95 95 86 95 MVRD
.MODEL MVRD NMOS VTO=-11.8 KP=24
LG 4 1 7N
.ENDS
*******
*SRC=BUZ-104;BUZ-104;MOSFETs N;Siemens;50V 17.5A 0.1 Ohm
*SYM=N-MOSFET
.SUBCKT BUZ-104 1 2 3
LS 5 2 7N
LD 97 3 5N
RG 95 96 7.4
RS 5 76 0.063
D104 76 97 DREV
.MODEL DREV D CJO=0.37N RS=20M TT=150N IS=300P BV=50
M104 98 96 76 76 MBUZ
.MODEL MBUZ NMOS VTO=3.5 KP=8.56
M2 96 98 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=.1
M3 98 96 8 8 MSW
COX 96 8 0.83N
DGD 8 98 DCGD
.MODEL DCGD D CJO=0.5N M=0.548 VJ=1.027
CGS 76 96 .36N
RD 98 97 0.004
LG 95 1 7N
.ENDS
*******
