*Aug 17, 2010
*Doc. ID: 90551, Rev. A
*File Name: irfz24ns_PS.txt and irfz24ns_PS.spi
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product datasheet.  Designers should refer to the
*appropriate data sheet of the same number for guaranteed specification
*limits.
.SUBCKT irfz24ns 1 2 3
* SPICE3 MODEL WITH THERMAL RC NETWORK
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Jul 17, 02
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.51818 LAMBDA=0 KP=6.23359
+CGSO=3e-06 CGDO=1e-07
RS 8 3 0.03
D1 3 1 MD
.MODEL MD D IS=2.13758e-11 RS=0.0118956 N=1.18924 BV=55
+IBV=0.00025 EG=1 XTI=2.43368 TT=0
+CJO=3e-10 VJ=1.73269 M=0.500012 FC=0.5
RDS 3 1 1e+06
RD 9 1 1e-05
RG 2 7 1.45002
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=4.19161e-10 VJ=0.5 M=0.59554 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 6.79024e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS irfz24ns

*SPICE Thermal Model Subcircuit
.SUBCKT irfz24nst 3 0
*(3 Layers)

R_RTHERM1         2 1  0.526
R_RTHERM2         3 2  1.048
R_RTHERM3         0 3  0.413
C_CTHERM1         1 0  0.000266
C_CTHERM2         0 2  0.00141
C_CTHERM3         3 0  0.050571

.ENDS irfz24nst


