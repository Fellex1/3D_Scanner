*IRF150 MCE 5/15/98
*100V  40A .045 ohm Power MOSFET pkg:TO-3 3,1,2
.SUBCKT IRF150   10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  20.4M
RS  40  3  2.12M
RG  20  2  3.75
CGS  2  3  1.65N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  4.49N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  12.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=208K THETA=60M ETA=2M VTO=3 KP=6.84)
.MODEL DCGD D (CJO=4.49N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=166N N=1.5 RS=43.8M BV=100 CJO=2.8N VJ=0.8 M=0.42 TT=600N)
.MODEL DLIM D (IS=100U)
.ENDS 


